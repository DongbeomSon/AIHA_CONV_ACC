`timescale 1ns / 1ps

module IFM_BUF (
    clk,
    stall,
    rst_n,
    ifm_input,
    ifm_read,
    ifm_buf0,
    ifm_buf1,
    ifm_buf2
);

    input clk;
    input stall;
    input rst_n;
    input signed [7:0] ifm_input;
    input ifm_read;
    output signed [7:0] ifm_buf0;
    output signed [7:0] ifm_buf1;
    output signed [7:0] ifm_buf2;

    reg signed [7:0] ifm_buf[2:0];

    integer i;

    always @(posedge clk or negedge rst_n)
        if (~rst_n) begin
            for (i = 0; i < 3; i = i + 1) begin
                ifm_buf[i] <= 0;
            end
        end else begin
            if (!stall) begin
                if (ifm_read) begin
                    ifm_buf[2] <= ifm_buf[1];
                    ifm_buf[1] <= ifm_buf[0];
                    ifm_buf[0] <= ifm_input;
                end else begin
                    ifm_buf[2] <= ifm_buf[2];
                    ifm_buf[1] <= ifm_buf[1];
                    ifm_buf[0] <= ifm_buf[0];
                end
            end
        end

    assign ifm_buf0 = ifm_buf[0];
    assign ifm_buf1 = ifm_buf[1];
    assign ifm_buf2 = ifm_buf[2];

endmodule
